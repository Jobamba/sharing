-- --------------------------------------------------------------------
--   $Id$ 
--   $Log$
--   Dateiname   : fir-a0-c0-cf.vhd
--   Titel       : Configuration fir_a0_c0 of fir ( a0 )
--   Ersteller   : dmpa
--   Projekt     : digitalmpa
--   Datum       : 27/11/19 13:14:03
--   Bemerkungen :
--               : $Log$
-- --------------------------------------------------------------------
-- library XXX ;

configuration fir_a1_c0 of fir is
  for a1

    -- Entity-Architecture Pairs Configurations
    -- for instance : component use entity work.entity(architecture) ;
    --    generic map(...) ;
    --    port map(...) ;
    -- end for ;

    -- Lower-Level Configurations
    -- for instance : component use configuration work.unit_con ;
    --    generic map(...) ;
    --    port map(...) ;
    -- end for ;

  end for ;
end fir_a1_c0;
